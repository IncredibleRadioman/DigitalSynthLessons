library IEEE; use IEEE.STD_LOGIC_1164.all;
use IEEE.STD_LOGIC_TEXTIO.ALL; use STD.TEXTIO.all;

entity testbench3 is
end;

architecture sim of testbench3 is
    component sillyfunction
    port(a, b, c: in STD_LOGIC;
        y: out STD_LOGIC);
    end component;

    signal a, b, c, y: STD_LOGIC;
    signal y_expected: STD_LOGIC;
    signal clk, reset: STD_LOGIC;
begin
    -- DUT
    dut: sillyfunction port map(a, b, c, y);
    -- generate clocks
    process begin
        clk <= '1'; wait for 5 ns;
        clk <= '0'; wait for 5 ns;
    end process;

    -- send reset after start
    process begin
        reset <= '1'; wait for 27 ns; reset <= '0';
        wait;
    end process;

    -- launch the test
    process is
        file tv: text;
        variable L: line;
        variable vector_in: std_logic_vector
            (2 downto 0);
        variable dummy: character;
        variable vector_out: std_logic;
        variable vectornum: integer := 0;
        variable errors: integer := 0;
    begin
        FILE_OPEN(tv, "example.tv", READ_MODE);
        while not endfile(tv) loop
            -- change vectors after posedge
            wait until rising_edge(clk);
            -- read the next string 
            readline(tv, L);
            read(L, vector_in);
            read(L, dummy);
            read(L, vector_out);
            (a, b, c) <= vector_in(2 downto 0)
                after 1 ns;
            y_expected <= vector_out after 1 ns;
            -- check results
            -- after negedge
            wait until falling_edge(clk);
            if y /= y_expected then
                report "Error: y = " & std_logic'image(y);
                errors := errors + 1;
            end if;
            vectornum := vectornum + 1;
        end loop;
        -- results
        if (errors = 0) then
            report "NO ERRORS -- " &
            integer'image(vectornum) &
            " tests completed successfully."
            severity failure;
        else
            report integer'image(vectornum) &
            " tests completed, errors = " &
            integer'image(errors)
            severity failure;
        end if;
    end process;
end;